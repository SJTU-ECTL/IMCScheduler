module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 ;
  assign n12 = x4 | x8 ;
  assign n13 = x1 & x4 ;
  assign n14 = n13 ^ x0 ^ 1'b0 ;
  assign n15 = ( x4 & ~n12 ) | ( x4 & n14 ) | ( ~n12 & n14 ) ;
  assign n16 = x6 | x7 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = x4 & x8 ;
  assign n19 = n17 | n18 ;
  assign n20 = ~x5 & n19 ;
  assign n21 = ( x3 & x4 ) | ( x3 & x7 ) | ( x4 & x7 ) ;
  assign n22 = x3 & ~x4 ;
  assign n23 = x1 & ~x2 ;
  assign n24 = x5 & ~x7 ;
  assign n25 = n23 & n24 ;
  assign n26 = x3 & ~n25 ;
  assign n27 = ( n21 & n22 ) | ( n21 & ~n26 ) | ( n22 & ~n26 ) ;
  assign n28 = ~x4 & x5 ;
  assign n29 = n27 ^ x8 ^ 1'b0 ;
  assign n30 = ( n27 & n28 ) | ( n27 & n29 ) | ( n28 & n29 ) ;
  assign n31 = n20 | n30 ;
  assign n32 = ~x9 & n31 ;
  assign n33 = x3 | x8 ;
  assign n34 = x7 ^ x4 ^ 1'b0 ;
  assign n35 = ( x7 & n33 ) | ( x7 & n34 ) | ( n33 & n34 ) ;
  assign n36 = n23 & ~n35 ;
  assign n37 = ~x1 & x2 ;
  assign n38 = x7 | x8 ;
  assign n39 = n37 & ~n38 ;
  assign n40 = x9 | n39 ;
  assign n41 = n36 | n40 ;
  assign n42 = ~x6 & n41 ;
  assign n43 = x6 & x9 ;
  assign n44 = n43 ^ x5 ^ 1'b0 ;
  assign n45 = ( n42 & n43 ) | ( n42 & n44 ) | ( n43 & n44 ) ;
  assign n46 = n32 | n45 ;
  assign n47 = ~x10 & n46 ;
  assign n48 = x3 ^ x2 ^ 1'b0 ;
  assign n49 = x8 | x9 ;
  assign n50 = n48 & ~n49 ;
  assign n51 = x10 | n50 ;
  assign n52 = ~x7 & n51 ;
  assign n53 = x9 & x10 ;
  assign n54 = x8 & n53 ;
  assign n55 = n52 | n54 ;
  assign n56 = x6 & n55 ;
  assign n57 = ~x6 & x10 ;
  assign n58 = x7 & n57 ;
  assign n59 = n56 | n58 ;
  assign n60 = n47 | n59 ;
  assign n61 = ( ~x2 & x4 ) | ( ~x2 & n49 ) | ( x4 & n49 ) ;
  assign n62 = ( x2 & x4 ) | ( x2 & ~n16 ) | ( x4 & ~n16 ) ;
  assign n63 = ~n61 & n62 ;
  assign n64 = x1 & n63 ;
  assign n65 = x4 & ~x8 ;
  assign n66 = x7 & ~x9 ;
  assign n67 = n65 & n66 ;
  assign n68 = n64 | n67 ;
  assign n69 = x3 & n68 ;
  assign n70 = x9 ^ x7 ^ 1'b0 ;
  assign n71 = ( x7 & n18 ) | ( x7 & ~n70 ) | ( n18 & ~n70 ) ;
  assign n72 = x6 & n71 ;
  assign n73 = n69 | n72 ;
  assign n74 = x8 & ~x9 ;
  assign n75 = n74 ^ n71 ^ x9 ;
  assign n76 = ~x6 & n75 ;
  assign n77 = ( x5 & n73 ) | ( x5 & n76 ) | ( n73 & n76 ) ;
  assign n78 = x4 | x9 ;
  assign n79 = x2 | x7 ;
  assign n80 = n78 & n79 ;
  assign n81 = x1 | n80 ;
  assign n82 = ( ~x0 & x2 ) | ( ~x0 & x7 ) | ( x2 & x7 ) ;
  assign n83 = x1 & x2 ;
  assign n84 = ( x0 & x7 ) | ( x0 & ~n83 ) | ( x7 & ~n83 ) ;
  assign n85 = n82 | n84 ;
  assign n86 = ( ~x4 & n81 ) | ( ~x4 & n85 ) | ( n81 & n85 ) ;
  assign n87 = ~n74 & n81 ;
  assign n88 = n86 & n87 ;
  assign n89 = x6 | n88 ;
  assign n90 = ( n33 & n49 ) | ( n33 & n78 ) | ( n49 & n78 ) ;
  assign n91 = ( x9 & n70 ) | ( x9 & ~n90 ) | ( n70 & ~n90 ) ;
  assign n92 = n89 & ~n91 ;
  assign n93 = ( x5 & ~n76 ) | ( x5 & n92 ) | ( ~n76 & n92 ) ;
  assign n94 = ~n77 & n93 ;
  assign n95 = x10 | n94 ;
  assign n96 = x6 & ~x9 ;
  assign n97 = ~x4 & n96 ;
  assign n98 = x5 & ~x6 ;
  assign n99 = ~x3 & n98 ;
  assign n100 = n97 | n99 ;
  assign n101 = ~x2 & n100 ;
  assign n102 = x4 & ~x6 ;
  assign n103 = x2 & x3 ;
  assign n104 = x4 & x6 ;
  assign n105 = n103 & n104 ;
  assign n106 = ( n96 & n102 ) | ( n96 & n105 ) | ( n102 & n105 ) ;
  assign n107 = x10 | n106 ;
  assign n108 = ~x1 & n98 ;
  assign n109 = ( ~x3 & n97 ) | ( ~x3 & n108 ) | ( n97 & n108 ) ;
  assign n110 = n107 | n109 ;
  assign n111 = n101 | n110 ;
  assign n112 = ~x7 & n111 ;
  assign n113 = n57 | n112 ;
  assign n114 = ~x8 & n113 ;
  assign n115 = x6 & x10 ;
  assign n116 = x7 & n115 ;
  assign n117 = n74 & n116 ;
  assign n118 = n114 | n117 ;
  assign n119 = n95 & ~n118 ;
  assign n120 = x0 & n102 ;
  assign n121 = n28 ^ x3 ^ 1'b0 ;
  assign n122 = ( n28 & n120 ) | ( n28 & ~n121 ) | ( n120 & ~n121 ) ;
  assign n123 = x1 & n122 ;
  assign n124 = x0 & x1 ;
  assign n125 = x3 & ~n124 ;
  assign n126 = x6 ^ x4 ^ 1'b0 ;
  assign n127 = ( x6 & ~n125 ) | ( x6 & n126 ) | ( ~n125 & n126 ) ;
  assign n128 = x5 | n127 ;
  assign n129 = ~n123 & n128 ;
  assign n130 = x2 & ~n129 ;
  assign n131 = x2 | x6 ;
  assign n132 = x5 ^ x3 ^ 1'b0 ;
  assign n133 = ( x5 & ~n131 ) | ( x5 & n132 ) | ( ~n131 & n132 ) ;
  assign n134 = x4 & n133 ;
  assign n135 = n130 | n134 ;
  assign n136 = ~x7 & n135 ;
  assign n137 = x3 & x4 ;
  assign n138 = ~x5 & x6 ;
  assign n139 = x2 & n138 ;
  assign n140 = n108 | n139 ;
  assign n141 = n137 & n140 ;
  assign n142 = x5 & x6 ;
  assign n143 = ~n137 & n142 ;
  assign n144 = n141 | n143 ;
  assign n145 = n136 | n144 ;
  assign n146 = ~x8 & n145 ;
  assign n147 = ~x6 & x7 ;
  assign n148 = x3 & n147 ;
  assign n149 = x6 & ~x7 ;
  assign n150 = ~x2 & n149 ;
  assign n151 = n148 | n150 ;
  assign n152 = x4 & x5 ;
  assign n153 = n151 & n152 ;
  assign n154 = x6 & x7 ;
  assign n155 = ~n152 & n154 ;
  assign n156 = n153 | n155 ;
  assign n157 = n146 | n156 ;
  assign n158 = ~x9 & n157 ;
  assign n159 = ( n24 & n104 ) | ( n24 & n147 ) | ( n104 & n147 ) ;
  assign n160 = ( x8 & n147 ) | ( x8 & n159 ) | ( n147 & n159 ) ;
  assign n161 = n158 | n160 ;
  assign n162 = ~x10 & n161 ;
  assign n163 = x5 & x9 ;
  assign n164 = x10 ^ x8 ^ 1'b0 ;
  assign n165 = ( x10 & n163 ) | ( x10 & ~n164 ) | ( n163 & ~n164 ) ;
  assign n166 = n154 & n165 ;
  assign n167 = x5 & x7 ;
  assign n168 = x8 & ~n167 ;
  assign n169 = x10 | n168 ;
  assign n170 = x9 & n169 ;
  assign n171 = n166 | n170 ;
  assign n172 = n162 | n171 ;
  assign n173 = ~x2 & n154 ;
  assign n174 = x5 & n18 ;
  assign n175 = n173 & n174 ;
  assign n176 = x5 | n12 ;
  assign n177 = n16 | n176 ;
  assign n178 = ~n175 & n177 ;
  assign n179 = x9 | x10 ;
  assign n180 = n178 | n179 ;
  assign n181 = x3 | n180 ;
  assign n182 = x5 | x6 ;
  assign n183 = n124 & ~n182 ;
  assign n184 = n159 | n183 ;
  assign n185 = n103 & n184 ;
  assign n186 = x7 & ~n142 ;
  assign n187 = ~n83 & n98 ;
  assign n188 = x9 | n187 ;
  assign n189 = n186 | n188 ;
  assign n190 = x4 | n149 ;
  assign n191 = ( ~x3 & x7 ) | ( ~x3 & n99 ) | ( x7 & n99 ) ;
  assign n192 = n190 & ~n191 ;
  assign n193 = ~n189 & n192 ;
  assign n194 = ~n185 & n193 ;
  assign n195 = x8 | n194 ;
  assign n196 = x7 & n142 ;
  assign n197 = ( ~x3 & x6 ) | ( ~x3 & x8 ) | ( x6 & x8 ) ;
  assign n198 = ( x2 & x3 ) | ( x2 & x6 ) | ( x3 & x6 ) ;
  assign n199 = n197 & n198 ;
  assign n200 = n167 & n199 ;
  assign n201 = x4 & n200 ;
  assign n202 = n196 ^ x9 ^ 1'b0 ;
  assign n203 = ( ~n196 & n201 ) | ( ~n196 & n202 ) | ( n201 & n202 ) ;
  assign n204 = n195 & ~n203 ;
  assign n205 = x10 | n204 ;
  assign n206 = x1 & x3 ;
  assign n207 = x0 & n206 ;
  assign n208 = x5 | x7 ;
  assign n209 = x8 | n208 ;
  assign n210 = n207 & ~n209 ;
  assign n211 = x8 & n167 ;
  assign n212 = ( n168 & n196 ) | ( n168 & n211 ) | ( n196 & n211 ) ;
  assign n213 = n210 | n212 ;
  assign n214 = x2 & n213 ;
  assign n215 = ( x3 & n99 ) | ( x3 & n212 ) | ( n99 & n212 ) ;
  assign n216 = n214 | n215 ;
  assign n217 = x4 & n216 ;
  assign n218 = ( n28 & n105 ) | ( n28 & n152 ) | ( n105 & n152 ) ;
  assign n219 = n218 ^ n98 ^ x6 ;
  assign n220 = ~n38 & n219 ;
  assign n221 = n179 | n220 ;
  assign n222 = n217 | n221 ;
  assign n223 = n179 | n218 ;
  assign n224 = n38 | n223 ;
  assign y0 = n60 ;
  assign y1 = n119 ;
  assign y2 = n172 ;
  assign y3 = n181 ;
  assign y4 = n205 ;
  assign y5 = n222 ;
  assign y6 = n224 ;
endmodule
